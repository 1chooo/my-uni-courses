LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SREGISTER IS
	PORT( SI, CK, CL : STD_LOGIC;
		  Q          : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END  SREGISTER;

ARCHITECTURE ARCH OF SREGISTER IS
BEGIN
	PROCESS(SI, CK, CL)
		VARIABLE REGT : STD_LOGIC_VECTOR(7 DOWNTO 0);
	BEGIN
		IF RISING_EDGE(CK) THEN
			IF CL = '1' THEN
				REGT := "00000000";
			ELSE
				REGT := REGT(6 DOWNTO 0) & SI;
			END IF;
			Q <= REGT;
		END IF;
	END PROCESS;
END ARCH;