LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE WORK.BIT_DEF.ALL;


ENTITY ACC IS
PORT (
		CLK     : IN  STD_LOGIC;
		RST     : IN  STD_LOGIC;
		RST_R   : IN  STD_LOGIC;
		S		: IN  STD_LOGIC;
		REG_IN  : IN  STD_LOGIC_VECTOR( DATA_WIDTH -1 DOWNTO 0);
		FINISH	: OUT STD_LOGIC;
		REG_OUT : OUT STD_LOGIC_VECTOR( DATA_WIDTH -1 DOWNTO 0);
	 );
END ACC;


ARCHITECTURE MIAT_REG_ARCH OF ACC IS
	SIGNAL REG : STD_LOGIC_VECTOR( DATA_WIDTH -1 DOWNTO 0);

BEGIN
	PROCESS(CLK)
	BEGIN
		IF RST = '0' OR RST_R = '1' THEN
			REG <= ( OTHERS => '0');
		ELSIF CLK'EVENT AND CLK = '1' THEN
			IF S = '1' THEN
				REG <= REG_IN;
				FINISH <= '1';
			END IF;
		END IF;
	END PROCESS;
	REG_OUT <= REG;
END MIAT_REG_ARCH;
