LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY BCDADDER IS
	PORT( A, B       : IN  INTEGER RANGE 0 TO 99;
		  Y2, Y1, Y0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END BCDADDER;

ARCHITECTURE ARCH OF BCDADDER IS
BEGIN
	PROCESS(A, B)
		VARIABLE SUM:INTEGER RANGE 0 TO 200;
		VARIABLE OUTPUT:STD_LOGIC_VECTOR(3 DOWNTO 0);
		VARIABLE TMP:INTEGER RANGE 0 TO 9;
	BEGIN
		SUM := A + B;
		TMP := SUM REM 10;
		DIG0 : FOR I IN 0 TO 3 LOOP
			IF ((TMP MOD 2) = 1) THEN OUTPUT(I) := '1';
			ELSE OUTPUT(I) := '0';
			END IF;
			TMP := TMP / 2;
		END LOOP;
		Y0 <= OUTPUT;
		
		TMP := (SUM / 10) REM 10;
		DIG1 : FOR I IN 0 TO 3 LOOP
			IF ((TMP MOD 2) = 1) THEN OUTPUT(I) := '1';
			ELSE OUTPUT(I) := '0';
			END IF;
			TMP := TMP/2;
		END LOOP;
		Y1 <= OUTPUT;
		
		TMP := (SUM / 100);
		DIG2: FOR I IN 0 TO 3 LOOP
			IF ((TMP MOD 2) = 1) THEN OUTPUT(I) := '1';
			ELSE OUTPUT(I) := '0';
			END IF;
			TMP := TMP / 2;
		END LOOP;
		Y2 <= OUTPUT;
	END PROCESS;
END ARCH;