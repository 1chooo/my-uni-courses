LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DEBOUNCING2 IS 
	PORT( DIN, CK : IN  STD_LOGIC;
			  DOUT    : OUT STD_LOGIC);
END DEBOUNCING2;

ARCHITECTURE ARCH OF DEBOUNCING2 IS
BEGIN
	PROCESS(CK)
		VARIABLE TMP : INTEGER RANGE 0 TO 9;
	BEGIN 
		IF RISING_EDGE(CK) THEN
		  IF DIN = '1' THEN
			   TMP := 0;
				 COUT <= '1';
			ELSE 
				TMP := TMP + 1;
				IF TMP = 4 THEN
					TMP := 0;
					DOUT <= '0';
				END IF;
			END IF;
		END IF;
	END PROCESS;
END ARCH;
