LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY COUNTER4B IS
	PORT(CL, PULSEIN : IN STD_LOGIC;
	     Q           : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END COUNTER4B;

ARCHITECTURE ARCH OF COUNTER4B IS
	COMPONENT DFF1
		PORT(CL, CK, T : IN STD_LOGIC;
		     Q , QBAR  : OUT STD_LOGIC);
	END COMPONENT;
	
	SIGNAL TMP : STD_LOGIC_VECTOR(4 DOWNTO 0);
	BEGIN
		TMP(0) <= PULSEIN;
		LP1 : FOR I IN 0 TO 3 GENERATE
			U : DFF1 PORT MAP (CL, TMP(I), '1', Q(I), TMP(I + 1));
		END GENERATE;
END ARCH;