LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MOD12 IS
	PORT( PULSEIN : IN STD_LOGIC;
		  Q       : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END MOD12;

ARCHITECTURE ARCH OF MOD12 IS
	COMPONENT DFF1
		PORT(CL, CK, T : IN STD_LOGIC;
		     Q , QBAR  : OUT STD_LOGIC);
	END COMPONENT;
	
	SIGNAL CL : STD_LOGIC;
	SIGNAL TMP1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
	SIGNAL TMP2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
	
BEGIN
	TMP1(0) <= PULSEIN;
	LP1 : FOR I IN 0 TO 3 GENERATE
		U : DFF1 PORT MAP (CL, TMP1(I), '1', TMP2(I), TMP1(I + 1));
	END GENERATE;
	CL <= TMP2(3) AND TMP2(2);
	Q <= TMP2;
END ARCH;