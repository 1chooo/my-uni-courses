LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ALU IS
PORT ( 
	  CLK, RST, S : IN  STD_LOGIC;
      A           : IN  STD_LOGIC;
      B           : IN  STD_LOGIC;
      F           : IN  STD_LOGIC_VECTOR( 3 DOWNTO 0 );
      O           : OUT STD_LOGIC
      );
END ALU;

ARCHITECTURE ACTION OF ALU IS
	SIGNAL REG : STD_LOGIC;

BEGIN 
	PROCESS(CLK)
	BEGIN
		IF RST = '0' THEN
			O <= '0';
		ELSIF CLK'EVENT AND CLK = '1' THEN
			IF S = '1' THEN
				0 <= REG;
			END IF;
		END IF;
	END PROCESS;

	REG <= NOT A  WHEN F = "0000" ELSE
	NOT (A OR B)  WHEN F = "0001" ELSE
	(NOT A) AND B WHEN F = "0010" ELSE 
	'0'           WHEN F = "0011" ELSE 
	NOT (A AND B) WHEN F = "0100" ELSE 
	NOT B         WHEN F = "0101" ELSE
	A XOR B       WHEN F = "0110" ELSE
	A AND (NOT B) WHEN F = "0111" ELSE
	(NOT A) OR B  WHEN F = "1000" ELSE
	NOT (A XOR B) WHEN F = "1001" ELSE
	B             WHEN F = "1010" ELSE
	A AND B       WHEN F = "1011" ELSE
	'1'           WHEN F = "1100" ELSE
	A OR (NOT B)  WHEN F = "1101" ELSE 
	A             WHEN F = "1111" ELSE
	'0';
END ACTION;
