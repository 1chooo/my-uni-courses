LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DEBOUNCING IS
  PORT( DIN, CK : IN  STD_LOGIC;
			  DOUT    : OUT STD_LOGIC);
END DEBOUNCING;

ARCHITECTURE ARCH OF DEBOUNCING IS
	COMPONENT DFF1
		PORT( D, CK : IN  STD_LOGIC;
				  Q     : OUT STD_LOGIC);
	END COMPONENT;

	SIGNAL TMP : STD_LOGIC_VECTOR(4 DOWNTO 0);
BEGIN
	TMP(0) <= DIN;
  LP1 : FOR I IN 1 TO 4 GENERATE
		 U1 : DFF1 PORT MAP(TMP(I - 1), CK, TMP(I));
	END GENERATE;

	DOUT <= TMP(4) AND TMP(3) AND TMP(2) AND TMP(1);
END ARCH;
