LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY MUX4TO1 IS
	PORT(
		A : IN  STD_LOGIC_VECTOR( 3 DOWNTO 0 );
		S : IN  STD_LOGIC_VECTOR( 1 DOWNTO 0 );
		Y : OUT STD_LOGIC
		);
END MUX4TO1;

ARCHITECTURE ARCH OF MUX4TO1 IS
BEGIN
	WITH S SELECT
	Y <= A(0) WHEN "00",
		  A(1) WHEN "01",
		  A(2) WHEN "10",
		  A(3) WHEN OTHERS;
END ARCH;